

`define SYNC_SIMPLE sync
`define SYNC_BLOCK  sync_block
`define SYNC_MERGE  sync_merge

// select one
`define MOD_SYNC `SYNC_BLOCK
