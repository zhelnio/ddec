
// select one
//`define SYNC_BLOCK
//`define SYNC_IMPL0
`define SYNC_IMPL1
